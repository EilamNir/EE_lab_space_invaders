// Design types
// =================

typedef logic signed [10:0] coordinate;
typedef logic signed [16:0] fixed_point; //TODO: Consider changing this to 16 bit, and changing FIXED_POINT_MULTIPLIER to 32 from 64
typedef logic [7:0] RGB;
typedef logic [28:0] VGA;
typedef logic [7:0] audio;
typedef logic [8:0] keycode;
typedef logic [6:0] hex_dig;
typedef logic [2:0] game_stage;
typedef logic [3:0] edge_code;
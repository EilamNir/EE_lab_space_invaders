//--------------------------------------
// (c) Technion IIT, Department of Electrical Engineering 2021 
//-- SystemVerilog version June 2018 Alex Grinshpun
// convert to 8 bits table - dudy march 2019 
//--------------------------------------


module	sintable	 #( 
					COUNT_SIZE = 8  // size of the table (in bits) 
		)	
		(	
//		--////////////////////	Clock Input	 	////////////////////	
					input		logic	clk,
					input		logic	resetN,
					input		logic [COUNT_SIZE-1:0]	addr,
					output	logic [15:0]	Q // table function output 
			);






localparam int table_size = (2**COUNT_SIZE)-1;

logic [7:0] tmp8bit  ; 

const logic [0:table_size-1] [7:0] sin_table = {

8'h00,
8'h06,
8'h0C,
8'h12,
8'h19,
8'h1F,
8'h25,
8'h2B,
8'h31,
8'h38,
8'h3E,
8'h44,
8'h4A,
8'h50,
8'h56,
8'h5C,
8'h61,
8'h67,
8'h6D,
8'h73,
8'h78,
8'h7E,
8'h83,
8'h88,
8'h8E,
8'h93,
8'h98,
8'h9D,
8'hA2,
8'hA7,
8'hAB,
8'hB0,
8'hB5,
8'hB9,
8'hBD,
8'hC1,
8'hC5,
8'hC9,
8'hCD,
8'hD1,
8'hD4,
8'hD8,
8'hDB,
8'hDE,
8'hE1,
8'hE4,
8'hE7,
8'hEA,
8'hEC,
8'hEE,
8'hF1,
8'hF3,
8'hF4,
8'hF6,
8'hF8,
8'hF9,
8'hFB,
8'hFC,
8'hFD,
8'hFE,
8'hFE,
8'hFF,
8'hFF,
8'hFF,
8'hFF,
8'hFF,
8'hFF,
8'hFF,
8'hFE,
8'hFE,
8'hFD,
8'hFC,
8'hFB,
8'hF9,
8'hF8,
8'hF6,
8'hF4,
8'hF3,
8'hF1,
8'hEE,
8'hEC,
8'hEA,
8'hE7,
8'hE4,
8'hE1,
8'hDE,
8'hDB,
8'hD8,
8'hD4,
8'hD1,
8'hCD,
8'hC9,
8'hC5,
8'hC1,
8'hBD,
8'hB9,
8'hB5,
8'hB0,
8'hAB,
8'hA7,
8'hA2,
8'h9D,
8'h98,
8'h93,
8'h8E,
8'h88,
8'h83,
8'h7E,
8'h78,
8'h73,
8'h6D,
8'h67,
8'h61,
8'h5C,
8'h56,
8'h50,
8'h4A,
8'h44,
8'h3E,
8'h38,
8'h31,
8'h2B,
8'h25,
8'h1F,
8'h19,
8'h12,
8'h0C,
8'h06,
8'h00,
8'hFA,
8'hF4,
8'hEE,
8'hE7,
8'hE1,
8'hDB,
8'hD5,
8'hCF,
8'hC8,
8'hC2,
8'hBC,
8'hB6,
8'hB0,
8'hAA,
8'hA4,
8'h9F,
8'h99,
8'h93,
8'h8D,
8'h88,
8'h82,
8'h7D,
8'h78,
8'h72,
8'h6D,
8'h68,
8'h63,
8'h5E,
8'h59,
8'h55,
8'h50,
8'h4B,
8'h47,
8'h43,
8'h3F,
8'h3B,
8'h37,
8'h33,
8'h2F,
8'h2C,
8'h28,
8'h25,
8'h22,
8'h1F,
8'h1C,
8'h19,
8'h16,
8'h14,
8'h12,
8'h0F,
8'h0D,
8'h0C,
8'h0A,
8'h08,
8'h07,
8'h05,
8'h04,
8'h03,
8'h02,
8'h02,
8'h01,
8'h01,
8'h01,
8'h00,
8'h01,
8'h01,
8'h01,
8'h02,
8'h02,
8'h03,
8'h04,
8'h05,
8'h07,
8'h08,
8'h0A,
8'h0C,
8'h0D,
8'h0F,
8'h12,
8'h14,
8'h16,
8'h19,
8'h1C,
8'h1F,
8'h22,
8'h25,
8'h28,
8'h2C,
8'h2F,
8'h33,
8'h37,
8'h3B,
8'h3F,
8'h43,
8'h47,
8'h4B,
8'h50,
8'h55,
8'h59,
8'h5E,
8'h63,
8'h68,
8'h6D,
8'h72,
8'h78,
8'h7D,
8'h82,
8'h88,
8'h8D,
8'h93,
8'h99,
8'h9F,
8'hA4,
8'hAA,
8'hB0,
8'hB6,
8'hBC,
8'hC2,
8'hC8,
8'hCF,
8'hD5,
8'hDB,
8'hE1,
8'hE7,
8'hEE,
8'hF4,
8'hFA
 };

 

always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN)
			tmp8bit	<= 8'h00;
	else 
		tmp8bit	<= sin_table[addr]; //  get sine (or other function) value from the table   

end

	assign 	Q = { {8{tmp8bit[7]}} ,  tmp8bit[7:0] }  ; // sign extend the msb  

endmodule

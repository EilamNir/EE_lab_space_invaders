module background
(
);

endmodule

// Design types
// =================

typedef logic signed [10:0] coordinate;
typedef logic [7:0] RGB;
module missiles
(
);

endmodule

module player
(
);

endmodule

module video_unit
(
);

endmodule

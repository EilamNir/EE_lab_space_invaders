module monsters
(
);

endmodule

module obstacles
(
);

endmodule

module sound_unit
(
);

endmodule

module hit_detection
(
);

endmodule

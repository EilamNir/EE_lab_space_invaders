// Design parameters
// =================

`include "types.sv"
